* SPICE 

V 3 0 DC 12

R0 1 0 100
R1 1 0 100
R3 2 1 100
R2 3 2 100
R4 3 2 100

.op
.tran 0 10ms 0ms 0.1ms
.print v(1) v(2) v(3) 
.end 
